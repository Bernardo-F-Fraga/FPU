module FPU (

input logic [31:0] a,
input logic [31:0] b,
input logic [1:0]  op,

output logic [31:0] res

);


endmodule